`ifndef VIP_RESET_PKG_SV
`define VIP_RESET_PKG_SV

package vip_reset_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "vip_reset_defines.sv"

    `include "vip_reset_types.sv"

    `include "seq/vip_reset_seq_item.sv"
    `include "seq/vip_reset_sequence.sv"

    `include "uvc/vip_reset_agent_configuration.sv"
    `include "uvc/vip_reset_monitor_item.sv"
    `include "uvc/vip_reset_monitor.sv"
    `include "uvc/vip_reset_driver.sv"
    `include "uvc/vip_reset_sequencer.sv"
    `include "uvc/vip_reset_agent.sv"

    `include "vip_reset_undefines.sv"
endpackage
`endif//VIP_RESET_PKG_SV