`ifndef VIP_RESET_UNDEFINES_SV
`define VIP_RESET_UNDEFINES_SV

`undef GETTER
`undef SETTER
`undef TESTER
`undef ACCESSOR
`undef GTN
`undef CHK
`undef CHK_FATAL
`undef CHK_RAND
`undef CHK_STD_RAND

`endif//VIP_RESET_UNDEFINES_SV